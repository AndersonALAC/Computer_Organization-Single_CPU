`timescale 1ns / 1ps

module ins_mem(
    input ins_addr,
    output [31:0] Inst_out
);


endmodule